package seq_pkg;
	import uvm_pkg::*;
	import ahb_pkg::*;
	import uart_pkg::*;

	`include"vip_tx_sequence.sv";
	`include"vip_tx_parity_error_sequence.sv";

endpackage

package env_pkg;

	import uvm_pkg::*;
	import apb_pkg::*;
	import axi_pkg::*;
	import bsc_regmodel_pkg::*;

	`include"scoreboard.sv";
	`include"environment.sv";
	`include"error_catcher.sv";

endpackage
